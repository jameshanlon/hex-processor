module processor
  (
    input logic i_rst,
    input logic i_clk
  );

endmodule
